// Copyright (c) 2023 - 2024 Meinhard Kissich
// SPDX-License-Identifier: MIT
// -----------------------------------------------------------------------------
// File  :  fazyrv_decode_mem1.sv
// Usage :  Instruction decoder optimized for 1 cycle memory delay.
//
// Param
//  - CHUNKSIZE       Data path width of the core.
//  - CONF            Configuration of the processor (MIN, INT, or CSR).
//  - RFTYPE          RAM type used for register file. Required in the control
//                    logic to adapt for delays.
//  - RST             Reduced reset type to save some more area.
//
// Ports
//  - clk_i               Clock input, sensitive to rising edge.
//  - rst_in              Reset, low active.
//  - trap_entry_i        Inform about trap.
//  - adr_lsbs_i          2 LSBs of the address for mask within a word.
//  - instr_i             Instruction word.
//  - stb_ir_i            Strobe instruction registers.
//  - stb_cntrl_i         Strobe control signals.
//  - cyc_two_i           In second operation cycle.
//  - shft_imm_i          Shift the immediate to the next CHUNKSIZE part.
//
//  - rs1_o               Address of source registers 1.
//  - rs2_o               Address of source registers 2.
//  - rd_o                Address of destination register.
//  - imm_o               CHUNKSIZE wide part of the immediate.
//
//  - alu_arith_o         ALU: arithmetic operation.
//  - alu_en_a_o          ALU: enable port a.
//  - alu_sub_o           ALU: arithmetical subtraction.
//  - alu_xor_o           ALU: logical xor.
//  - alu_and_o           ALU: logical and.
//  - alu_cmp_sign_o      ALU: consider sign bit for comparisons.
//  - alu_cmp_eq_o        ALU: if comparison, then check for equality.
//  - alu_cmp_inv_o       ALU: invert the comparison result.
//
//  - alu_aux_rev_o       ALU: reverse the ALU inputs.
//  - alu_aux_rs_a_pc_o   ALU: input the PC at input a, otherwise rs1.
//  - alu_aux_rs_b_imm_o  ALU: input the immediate at the a input,
//                        otherwise rs2.
//  - alu_aux_b_spm_d_o   ALU: input the spm_d output at the b input (has prio).
//  - alu_aux_use_cmp_o   ALU: use the comparison result as the output.
//
//  - ls_mask_o           Load and store mask.
//  - ld_sext_o           Sign-extend loaded data.
//  - sext_o              Inform spm_d to sign extend the data.
//
//  - rf_we_o             Rd in register file shall be written.
//
//  - instr_ld_o          Is load instruction.
//  - instr_st_o          Is store instruction.
//  - ls_b_o              If load or store, then we consider a byte.
//  - ls_h_o              If load or store, then we consider a half-word.
//  - ls_w_o              If load or store, then we consider a word.
//  - instr_shft_o        Is shift instruction.
//  - instr_left_o        Shift left in the spm_d.
//  - instr_any_br_o      Is a branch instruction.
//  - instr_jmp_o         Is a jump instruction.
//  - instr_slt_o         Is a set less than instruction.
//  - instr_csr_o         Is an isntruction that modifes a CSR.
//
//  - csr_hpmtc_o         Select hpm or timer counter instead of RF CSRs.
//  - csr_6_o             Write to a CSR with 6th CSR bit high.
//  - csr_high_o          Read high part of 64-bit hpmtc.
//
//  - mret_o              Is return from trap.
//  - mcause30_o          mcause part generated by decoder.
//  - except_o            Illegal instruction and/or ecall/ebreak
//                        (may be ignored, depending on CONF).
// -----------------------------------------------------------------------------

module fazyrv_decode_mem1 #(
  parameter CHUNKSIZE = 2,
  parameter CONF      = "MIN",
  parameter RFTYPE    = "BRAM_DP_BP",
  parameter RST       = "MIN"
) (
  input  logic              clk_i,
  input  logic              rst_in,
  input  logic              trap_entry_i,
  input  logic [1:0]        adr_lsbs_i,
  input  logic [31:0]       instr_i,
  input  logic              stb_ir_i,
  input  logic              stb_cntrl_i,
  input  logic              cyc_two_i,
  input  logic              shft_imm_i,

  output logic [4:0]            rs1_o,
  output logic [4:0]            rs2_o,
  output logic [4:0]            rd_o,
  output logic [CHUNKSIZE-1:0]  imm_o,

  output logic              alu_arith_o,
  output logic              alu_en_a_o,
  output logic              alu_sub_o,
  output logic              alu_xor_o,
  output logic              alu_and_o,
  output logic              alu_cmp_sign_o,
  output logic              alu_cmp_eq_o,
  output logic              alu_cmp_inv_o,

  output logic              alu_aux_rev_o,
  output logic              alu_aux_rs_a_pc_o,
  output logic              alu_aux_rs_b_imm_o,
  output logic              alu_aux_b_spm_d_o,
  output logic              alu_aux_use_cmp_o,

  output logic [3:0]        ls_mask_o,
  output logic              ld_sext_o,
  output logic              sext_o,

  output logic              rf_we_o,

  output logic              instr_ld_o,
  output logic              instr_st_o,
  output logic              ls_b_o,
  output logic              ls_h_o,
  output logic              ls_w_o,
  output logic              instr_shft_o,
  output logic              instr_left_o,
  output logic              instr_any_br_o,
  output logic              instr_jmp_o,
  output logic              instr_slt_o,
  output logic              instr_csr_o,

  output logic              csr_hpmtc_o,
  output logic              csr_6_o,
  output logic              csr_high_o,

  output logic              mret_o,
  output logic [1:0]        mcause30_o,
  output logic              except_o
);

// If 1, a smaller decoder is implemented. However, this
// leads to a reduced fmax
localparam SMALL = 1;

// --- misc ---

logic in_cycle_2;
assign in_cycle_2 = cyc_two_i;

// --- register decoding ---

logic [4:0] rs1_r;
logic [4:0] rs2_r;
logic [4:0] rd_r;

always_ff @(posedge clk_i) begin
  if (~rst_in & (RST != "MIN")) begin
    rs1_r <= 'b0;
    rs2_r <= 'b0;
    rd_r  <= 'b0;
  end else if (stb_ir_i) begin
    rs1_r <= instr_i[19:15];
    rs2_r <= instr_i[24:20];
    rd_r  <= instr_i[11:7];
  end
end

assign rs1_o = stb_ir_i ? instr_i[19:15] : rs1_r;
assign rs2_o = stb_ir_i ? instr_i[24:20] : rs2_r;
assign rd_o  = stb_ir_i ? instr_i[11:7]  : rd_r;

// --- imm decoding ---

logic [31:0] imm_r, imm_n;

logic [31:0] u_imm;
logic [31:0] j_imm;
logic [31:0] i_imm;
logic [31:0] s_imm;
logic [31:0] b_imm;

assign i_imm = { {21{instr_i[31]}}, instr_i[30:20] };
assign s_imm = { {21{instr_i[31]}}, instr_i[30:25], instr_i[11:7] };
assign b_imm = { {20{instr_i[31]}}, instr_i[7], instr_i[30:25],
                  instr_i[11:8], 1'd0};
assign u_imm = { instr_i[31:12], 12'd0 };
assign j_imm = { {12{instr_i[31]}}, instr_i[19:12], instr_i[20],
                  instr_i[30:21], 1'd0 };

logic is_u_imm;
logic is_j_imm;
logic is_i_imm;
logic is_s_imm;
logic is_b_imm;

// TODO: MRET compare are with passthrough + nop in current insn to use
// inc(pc) instead of alu to increment

/* svlint off style_keyword_1or2space */
/* svlint off style_keyword_construct */
/* svlint off style_keyword_1space */
always_comb begin
  imm_n = 32'd4;
  if (is_u_imm) imm_n = u_imm;
  else if (is_j_imm) imm_n = j_imm;
  else if (is_i_imm) imm_n = i_imm;
  else if (is_s_imm) imm_n = s_imm;
  else if (is_b_imm) imm_n = b_imm;
end
/* svlint on style_keyword_1or2space */
/* svlint on style_keyword_construct */
/* svlint on style_keyword_1space */


always_ff @(posedge clk_i) begin
  if (stb_ir_i) begin
    imm_r <= imm_n;
  end else if (shft_imm_i) begin
    imm_r <= {{CHUNKSIZE{1'bx}}, imm_r[31:CHUNKSIZE]};
  end
end

assign imm_o = imm_r[CHUNKSIZE-1:0];

// --- masks ---

always_ff @(posedge clk_i) begin
  if (stb_ir_i) begin
    ls_w_o    <= instr_i[13];
    ls_h_o    <= instr_i[12];
    ls_b_o    <= ~instr_i[13] & ~instr_i[12];

    ld_sext_o <= instr_i[14];
    sext_o    <= (~instr_i[14] & ~instr_i[4]) | (instr_i[30] & instr_i[4]);
  end
end

// Smaller than version below, inspired by SERV
assign ls_mask_o[3] = (adr_lsbs_i == 2'b11) | ls_w_o | (ls_h_o & adr_lsbs_i[1]);
assign ls_mask_o[2] = (adr_lsbs_i == 2'b10) | ls_w_o;
assign ls_mask_o[1] = (adr_lsbs_i == 2'b01) | ls_w_o | (ls_h_o & !adr_lsbs_i[1]);
assign ls_mask_o[0] = (adr_lsbs_i == 2'b00);


generate
  if (SMALL) begin
    always_comb begin
      is_b_imm = 1'b0;
      is_s_imm = 1'b0;
      is_i_imm = 1'b0;
      is_j_imm = 1'b0;
      is_u_imm = 1'b0;

      if (instr_i[2] & instr_i[3])
        is_j_imm = 1'b1;
      else if (~instr_i[2] & ~instr_i[4] & instr_i[6])
        is_b_imm = 1'b1;
      else if (instr_i[2] & ~instr_i[6])
        is_u_imm = 1'b1;
      else if (~instr_i[2] & ~instr_i[4] & instr_i[5])
        is_s_imm = 1'b1;
      // This does not work for csrrxi anymore, but fixes mret efficiently
      //else if (~(instr_i[4] & instr_i[5] & ~instr_i[6]))
      else if (~(instr_i[4] & instr_i[5]))
        is_i_imm = 1'b1;

    end
  end else begin

    assign is_b_imm = (!instr_i[13]&instr_i[6]&instr_i[5]&!instr_i[4]&
        !instr_i[3]&!instr_i[2]&instr_i[1]&instr_i[0]) | (
        instr_i[14]&instr_i[6]&instr_i[5]&!instr_i[4]&!instr_i[3]
        &!instr_i[2]&instr_i[1]&instr_i[0]);

    assign is_s_imm = (!instr_i[14]&!instr_i[12]&!instr_i[6]&instr_i[5]&
        !instr_i[4]&!instr_i[3]&!instr_i[2]
        &instr_i[1]&instr_i[0]) | (!instr_i[14]&!instr_i[13]&!instr_i[6]&
        instr_i[5]&!instr_i[4]&!instr_i[3]
        &!instr_i[2]&instr_i[1]&instr_i[0]);

    assign is_i_imm = (!instr_i[31]&!instr_i[30]&!instr_i[29]&!instr_i[28]&
    !instr_i[27]&!instr_i[26]&!instr_i[25]&!instr_i[6]&!instr_i[5]&instr_i[4
    ]&!instr_i[3]&!instr_i[2]&instr_i[1]&instr_i[0]) | (!instr_i[31]
        &!instr_i[29]&!instr_i[28]&!instr_i[27]&!instr_i[26]&!instr_i[25]&
        instr_i[14]&!instr_i[6]&!instr_i[5]
        &instr_i[4]&!instr_i[3]&!instr_i[2]&instr_i[1]&instr_i[0]) |
        (!instr_i[12]&!instr_i[6]&!instr_i[5]
        &instr_i[4]&!instr_i[3]&!instr_i[2]&instr_i[1]&instr_i[0]) |
        (!instr_i[14]&!instr_i[13]&!instr_i[12]
        &instr_i[6]&instr_i[5]&!instr_i[4]&!instr_i[3]&instr_i[2]&
        instr_i[1]&instr_i[0]) | (!instr_i[14]
        &!instr_i[12]&!instr_i[6]&!instr_i[5]&!instr_i[3]&!instr_i[2]&
        instr_i[1]&instr_i[0]) | (!instr_i[13]
        &!instr_i[6]&!instr_i[5]&!instr_i[4]&!instr_i[3]&!instr_i[2]&
        instr_i[1]&instr_i[0]) | (instr_i[13]
        &!instr_i[6]&!instr_i[5]&instr_i[4]&!instr_i[3]&!instr_i[2]&
        instr_i[1]&instr_i[0]);

    assign is_j_imm = (instr_i[6]&instr_i[5]&!instr_i[4]&instr_i[3]&
    instr_i[2]&instr_i[1]&instr_i[0]);

    assign is_u_imm = (!instr_i[6]&instr_i[4]&!instr_i[3]&instr_i[2]&
    instr_i[1]&instr_i[0]);
end
endgenerate

// --- store opcode ---

// Let the tool optimize away the bits that are not needed
logic [31:0] i_r;

always_ff @(posedge clk_i) begin
  if (~rst_in) begin
    // either to instr_i or to NOP, all 0s causes trap
    i_r <= instr_i; // 'b0;
  end else if (stb_ir_i) begin
    i_r <= instr_i;
  end
end

logic [31:0] ins;
logic stb_cntrl;

generate
  /* verilator lint_off WIDTHEXPAND */
  if (RFTYPE == "BRAM_DP_BP") begin
  /* verilator lint_on WIDTHEXPAND */
    assign ins = stb_ir_i ? instr_i : i_r;
    assign stb_cntrl = stb_cntrl_i | stb_ir_i;
  end else begin
    assign ins = i_r;
    assign stb_cntrl = stb_cntrl_i;
  end
endgenerate


always_ff @(posedge clk_i) begin
  if (stb_cntrl) begin
  alu_aux_b_spm_d_o <= (!ins[14]&!ins[12]&!ins[6]&!ins[5]&!ins[4]&in_cycle_2) | (
      !trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]&!ins[2]
      &in_cycle_2) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&!ins[5]&ins[4]
      &!ins[3]&!ins[2]) | (!trap_entry_i&!ins[13]&!ins[6]&!ins[5]&!ins[4]
      &in_cycle_2);

  alu_aux_rs_b_imm_o <= (!trap_entry_i&ins[13]&ins[12]&!ins[6]&!ins[5]
      &ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&ins[29]&!ins[14]&!ins[13]
      &!ins[12]&ins[6]&ins[4]) | (ins[14]&ins[6]&!ins[4]&!ins[3]&in_cycle_2) | (
      !ins[13]&ins[6]&!ins[4]&!ins[3]&in_cycle_2) | (!trap_entry_i&!ins[14]
      &!ins[12]&!ins[6]&!ins[4]&!in_cycle_2) | (!trap_entry_i&!ins[12]
      &!ins[6]&!ins[5]&ins[4]&!ins[3]&!ins[2]) | (!ins[13]&!ins[6]&!ins[5]
      &!ins[3]&!in_cycle_2) | (!trap_entry_i&!ins[14]&!ins[13]&!ins[6]
      &!ins[4]&!in_cycle_2) | (!trap_entry_i&ins[6]&!ins[4]&ins[2]
      &!in_cycle_2) | (!trap_entry_i&!ins[13]&!ins[6]&!ins[5]&!ins[4]
      &!in_cycle_2) | (!trap_entry_i&!ins[6]&!ins[5]&ins[4]&!ins[3]&ins[2]) | (
      !ins[6]&ins[5]&ins[4]&ins[2]);

  alu_aux_rs_a_pc_o <= (ins[14]&ins[6]&!ins[4]&!ins[3]&in_cycle_2) | (
      !ins[13]&ins[6]&!ins[4]&!ins[3]&in_cycle_2) | (!trap_entry_i&ins[6]
      &!ins[4]&ins[3]&ins[2]) | (ins[6]&!ins[4]&ins[2]&in_cycle_2) | (
      !trap_entry_i&!ins[6]&!ins[5]&ins[4]&!ins[3]&ins[2]) | (trap_entry_i);

  alu_aux_rev_o <= (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]
      &!ins[2]&!in_cycle_2) | (!ins[13]&!ins[6]&!ins[5]&!ins[3]&!in_cycle_2) | (
      !ins[14]&ins[6]&ins[4]&!in_cycle_2) | (ins[6]&!ins[4]&ins[2]
      &in_cycle_2) | (trap_entry_i);

  alu_cmp_inv_o <= (ins[14]&ins[12]&ins[6]&!ins[4]&!ins[3]) | (!ins[14]
      &!ins[13]&ins[12]&!ins[3]);

  alu_cmp_eq_o <= (!ins[14]&!ins[13]&!ins[3]);

  alu_cmp_sign_o <= (!trap_entry_i&!ins[12]&!ins[6]&!ins[5]&ins[4]&!ins[3]
      &!ins[2]) | (!trap_entry_i&!ins[12]&!ins[6]&ins[5]&ins[4]&!ins[2]) | (
      !trap_entry_i&!ins[13]&ins[6]&!ins[4]&!ins[3]&!ins[2]);

  alu_and_o <= (!trap_entry_i&ins[13]&ins[12]&!ins[6]&!ins[5]&ins[4]&!ins[3]
      &!ins[2]) | (!trap_entry_i&ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]
      &!ins[2]);

  alu_xor_o <= (!trap_entry_i&!ins[13]&!ins[6]&ins[5]&ins[4]) | (
      !trap_entry_i&!ins[13]&!ins[6]&ins[4]&!ins[3]);

  alu_sub_o <= (!trap_entry_i&ins[30]&!ins[12]&!ins[6]&ins[5]&ins[4]&!ins[2]);

  alu_en_a_o <= (!trap_entry_i&ins[13]&ins[12]&!ins[6]&!ins[5]&ins[4]&!ins[3]
      &!ins[2]) | (!trap_entry_i&ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]
      &!ins[2]) | (!trap_entry_i&ins[29]&!ins[14]&!ins[13]&!ins[12]&ins[6]
      &ins[4]) | (!trap_entry_i&!ins[14]&!ins[12]&!ins[6]&!ins[4]
      &!in_cycle_2) | (!trap_entry_i&ins[14]&ins[6]&!ins[4]&!ins[3]&!ins[2]) | (
      !trap_entry_i&!ins[12]&!ins[6]&!ins[5]&ins[4]&!ins[3]&!ins[2]) | (
      !trap_entry_i&!ins[14]&!ins[13]&!ins[6]&!ins[4]&!in_cycle_2) | (
      !trap_entry_i&!ins[12]&!ins[6]&ins[5]&ins[4]&!ins[2]) | (
      !trap_entry_i&ins[6]&!ins[4]&ins[2]&!in_cycle_2) | (!trap_entry_i
      &!ins[13]&ins[6]&!ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&!ins[13]
      &!ins[6]&!ins[5]&!ins[4]&!in_cycle_2) | (!trap_entry_i&!ins[6]&!ins[5]
      &ins[4]&!ins[3]&ins[2]);

  alu_arith_o <= (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]
      &!ins[2]&in_cycle_2) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]
      &ins[4]&!ins[2]&!in_cycle_2) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]
      &!ins[5]&ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&ins[29]&!ins[14]
      &!ins[13]&!ins[12]&ins[6]&ins[4]) | (!trap_entry_i&ins[14]&ins[6]
      &!ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&!ins[14]&!ins[12]&!ins[6]
      &ins[5]&!ins[4]) | (!trap_entry_i&ins[6]&!ins[4]&ins[3]&ins[2]) | (
      !trap_entry_i&!ins[14]&!ins[13]&!ins[6]&ins[5]&!ins[4]) | (
      !trap_entry_i&!ins[13]&ins[6]&!ins[4]&!ins[3]&!ins[2]) | (
      !trap_entry_i&!ins[14]&!ins[12]&!ins[6]&!ins[5]&!ins[4]) | (
      !trap_entry_i&!ins[13]&!ins[6]&!ins[5]&!ins[4]&in_cycle_2) | (
      !trap_entry_i&ins[6]&!ins[4]&!ins[3]&ins[2]) | (!trap_entry_i&!ins[13]
      &!ins[6]&!ins[5]&!ins[4]&!in_cycle_2) | (!trap_entry_i&!ins[14]
      &ins[13]&ins[6]&ins[4]) | (!trap_entry_i&!ins[14]&!ins[6]&ins[5]
      &ins[4]) | (!trap_entry_i&!ins[14]&ins[12]&ins[6]&ins[4]) | (
      !trap_entry_i&!ins[14]&!ins[6]&ins[4]&!ins[3]) | (!trap_entry_i
      &!ins[6]&!ins[5]&ins[4]&!ins[3]&ins[2]) | (!ins[6]&ins[5]&ins[4]
      &ins[2]) | (trap_entry_i);

  instr_jmp_o <= (!trap_entry_i&ins[6]&!ins[4]&ins[3]&ins[2]) | (
      !trap_entry_i&ins[6]&!ins[4]&!ins[3]&ins[2]);

  instr_any_br_o <= (!trap_entry_i&ins[14]&ins[6]&!ins[4]&!ins[3]&!ins[2]) | (
      !trap_entry_i&!ins[13]&ins[6]&!ins[4]&!ins[3]&!ins[2]);

  alu_aux_use_cmp_o <= (!trap_entry_i&!ins[14]&ins[13]&!ins[6]&ins[5]&ins[4]
      &!ins[2]) | (!trap_entry_i&!ins[14]&ins[13]&!ins[6]&ins[4]&!ins[3]
      &!ins[2]);

  instr_left_o <= (!trap_entry_i&!ins[14]&!ins[6]&ins[5]&ins[4]) | (
      !trap_entry_i&!ins[14]&!ins[6]&ins[4]&!ins[3]);

  instr_shft_o <= (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]
      &!ins[2]&in_cycle_2) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]
      &ins[4]&!ins[2]&!in_cycle_2) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]
      &!ins[5]&ins[4]&!ins[3]&!ins[2]);

  instr_st_o <= (!trap_entry_i&!ins[14]&!ins[12]&!ins[6]&ins[5]&!ins[4]) | (
      !trap_entry_i&!ins[14]&!ins[13]&!ins[6]&ins[5]&!ins[4]);

  instr_ld_o <= (!trap_entry_i&!ins[14]&!ins[12]&!ins[6]&!ins[5]&!ins[4]) | (
      !trap_entry_i&!ins[13]&!ins[6]&!ins[5]&!ins[4]&in_cycle_2) | (
      !trap_entry_i&!ins[13]&!ins[6]&!ins[5]&!ins[4]&!in_cycle_2);

  instr_slt_o <= (!trap_entry_i&!ins[14]&ins[13]&!ins[6]&ins[5]&ins[4]
      &!ins[2]) | (!trap_entry_i&!ins[14]&ins[13]&!ins[6]&ins[4]&!ins[3]
      &!ins[2]);

  rf_we_o <= (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]&!ins[2]
      &in_cycle_2) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]&ins[5]&ins[4]
      &!ins[2]&!in_cycle_2) | (!trap_entry_i&ins[13]&ins[12]&!ins[6]&!ins[5]
      &ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&ins[13]&ins[12]&!ins[6]
      &ins[5]&ins[4]&!ins[2]) | (!trap_entry_i&!ins[13]&ins[12]&!ins[6]
      &!ins[5]&ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&!ins[12]&!ins[6]
      &!ins[5]&ins[4]&!ins[3]&!ins[2]) | (!trap_entry_i&!ins[12]&!ins[6]
      &ins[5]&ins[4]&!ins[2]) | (ins[6]&!ins[4]&ins[2]&in_cycle_2) | (
      !trap_entry_i&!ins[14]&!ins[12]&!ins[6]&!ins[5]&!ins[4]) | (
      !trap_entry_i&!ins[13]&!ins[6]&!ins[5]&!ins[4]&in_cycle_2) | (
      !trap_entry_i&!ins[14]&ins[13]&ins[6]&ins[4]) | (!trap_entry_i
      &!ins[14]&ins[12]&ins[6]&ins[4]) | (!trap_entry_i&!ins[6]&!ins[5]
      &ins[4]&!ins[3]&ins[2]) | (!ins[6]&ins[5]&ins[4]&ins[2]) | (
      trap_entry_i);
  end
end

generate
  if (CONF == "CSR") begin
    always_ff @(posedge clk_i) begin
      instr_csr_o <= (!trap_entry_i&!ins[14]&ins[13]&ins[6]&ins[5]&ins[4]&!ins[3]
      &!ins[2]) | (!trap_entry_i&!ins[14]&ins[12]&ins[6]&ins[5]&ins[4]
      &!ins[3]&!ins[2]);
    end
    assign csr_hpmtc_o  = ins[31];
    assign csr_6_o      = ins[26];
    assign csr_high_o   = ins[27];
  end else begin
    assign instr_csr_o  = 1'b0;
    assign csr_hpmtc_o  = 1'b0;
    assign csr_6_o      = 1'b0;
    assign csr_high_o   = 1'b0;
  end

  if ((CONF == "INT") | (CONF == "CSR")) begin
    always_ff @(posedge clk_i) begin
      mret_o <= (!trap_entry_i&ins[29]&!ins[14]&!ins[13]&!ins[12]&ins[6]&ins[4]);
    end
  end else begin
    assign mret_o = 1'b0;
  end
endgenerate

// --- csr and trap ---

generate
  if ((CONF == "CSR") || (CONF == "INT")) begin
    // Illegal instruction: all 0s or all 1s, others might fail to be detected
    // due to area optimization.
    logic trap_insn;
    logic trap_e;

    always_ff @(posedge clk_i) begin
      trap_insn     <= (&ins[6:3]) | ~(|ins[1:0]);
      trap_e        <= (&ins[6:4]) &  ~(|ins[14:12]) & ~ins[29];
      mcause30_o[1] <= (&ins[6:4]) &  ~(|ins[14:12]) & ~ins[29] & ins[20];
      mcause30_o[0] <= (&ins[6:4]) &  ~(|ins[14:12]) & ~ins[29];
    end
    assign except_o   = trap_insn | trap_e;

    // 2  0010 ... illegal instr
    // 3  0011 ... break
    // 11 1011 ... ecall

  end else begin
    assign except_o     = 1'b0;
    assign mcause30_o   = 2'b0;
  end
endgenerate


endmodule
