// Copyright (c) 2023 - 2024 Meinhard Kissich
// SPDX-License-Identifier: MIT
// -----------------------------------------------------------------------------
// File  :  fazyrv_decode.sv
// Usage :  Instruction decoder.
//
// Param
//  - CHUNKSIZE       Data path width of the core.
//  - CONF            Configuration of the processor (MIN, INT, or CSR).
//  - RFTYPE          RAM type used for register file. Required in the control
//                    logic to adapt for delays.
//  - RST             Reduced reset type to save some more area. 
//
// Ports
//  - clk_i               Clock input, sensitive to rising edge.
//  - rst_in              Reset, low active.
//  - trap_entry_i        Inform about trap.
//  - adr_lsbs_i          2 LSBs of the address for mask within a word.
//  - instr_i             Instruction word.
//  - stb_ir_i            Strobe instruction registers.
//  - stb_cntrl_i         Strobe control signals.
//  - cyc_two_i           In second operation cycle.
//  - shft_imm_i          Shift the immediate to the next CHUNKSIZE part.
//
//  - rs1_o               Address of source registers 1.
//  - rs2_o               Address of source registers 2.
//  - rd_o                Address of destination register.
//  - imm_o               CHUNKSIZE wide part of the immediate.
//
//  - alu_arith_o         ALU: arithmetic operation.
//  - alu_en_a_o          ALU: enable port a.
//  - alu_sub_o           ALU: arithmetical subtraction.
//  - alu_xor_o           ALU: logical xor.
//  - alu_and_o           ALU: logical and.
//  - alu_cmp_sign_o      ALU: consider sign bit for comparisons.
//  - alu_cmp_eq_o        ALU: if comparison, then check for equality.
//  - alu_cmp_inv_o       ALU: invert the comparison result.
//
//  - alu_aux_rev_o       ALU: reverse the ALU inputs.
//  - alu_aux_rs_a_pc_o   ALU: input the PC at input a, otherwise rs1.
//  - alu_aux_rs_b_imm_o  ALU: input the immediate at the a input,
//                        otherwise rs2.
//  - alu_aux_b_spm_d_o   ALU: input the spm_d output at the b input (has prio).
//  - alu_aux_use_cmp_o   ALU: use the comparison result as the output.
//
//  - ls_mask_o           Load and store mask.
//  - ld_sext_o           Sign-extend loaded data.
//  - sext_o              Inform spm_d to sign extend the data.
//
//  - rf_we_o             Rd in register file shall be written.
//
//  - instr_ld_o          Is load instruction.
//  - instr_st_o          Is store instruction.
//  - ls_b_o              If load or store, then we consider a byte.
//  - ls_h_o              If load or store, then we consider a half-word.
//  - ls_w_o              If load or store, then we consider a word.
//  - instr_shft_o        Is shift instruction.
//  - instr_left_o        Shift left in the spm_d.
//  - instr_any_br_o      Is a branch instruction.
//  - instr_jmp_o         Is a jump instruction.
//  - instr_slt_o         Is a set less than instruction.
//  - instr_csr_o         Is an isntruction that modifes a CSR.
//  - ccx_o               Is chunked custom instruction.
//  - ccx_sel_o           Select custom instructions (part of func3).
//
//  - csr_hpmtc_o         Select hpm or timer counter instead of RF CSRs.
//  - csr_6_o             Write to a CSR with 6th CSR bit high.
//  - csr_high_o          Read high part of 64-bit hpmtc.
//
//  - mret_o              Is return from trap.
//  - mcause30_o          mcause part generated by decoder.
//  - except_o            Illegal instruction and/or ecall/ebreak
//                        (may be ignored, depending on CONF).

module fazyrv_decode #(
  parameter CHUNKSIZE = 2,
  parameter CONF = "MIN",
  parameter RST = "MIN"
) (
  input  logic              clk_i,
  input  logic              rst_in,
  input  logic              trap_entry_i,
  input  logic [1:0]        adr_lsbs_i,
  input  logic [31:0]       instr_i,
  input  logic              stb_ir_i,
  input  logic              stb_cntrl_i,
  input  logic              cyc_two_i,
  input  logic              shft_imm_i,

  output logic [4:0]            rs1_o,
  output logic [4:0]            rs2_o,
  output logic [4:0]            rd_o,
  output logic [CHUNKSIZE-1:0]  imm_o,

  output logic              alu_arith_o,
  output logic              alu_en_a_o,
  output logic              alu_sub_o,
  output logic              alu_xor_o,
  output logic              alu_and_o,
  output logic              alu_cmp_sign_o,
  output logic              alu_cmp_eq_o,
  output logic              alu_cmp_inv_o,

  output logic              alu_aux_rev_o,
  output logic              alu_aux_rs_a_pc_o,
  output logic              alu_aux_rs_b_imm_o,
  output logic              alu_aux_b_spm_d_o,
  output logic              alu_aux_use_cmp_o,

  output logic [3:0]        ls_mask_o,
  output logic              ld_sext_o,
  output logic              sext_o,

  output logic              rf_we_o,

  output logic              instr_ld_o,
  output logic              instr_st_o,
  output logic              ls_b_o,
  output logic              ls_h_o,
  output logic              ls_w_o,
  output logic              instr_shft_o,
  output logic              instr_left_o,
  output logic              instr_any_br_o,
  output logic              instr_jmp_o,
  output logic              instr_slt_o,
  output logic              instr_csr_o,

  output logic              ccx_o,
  output logic [1:0]        ccx_sel_o,

  output logic              csr_hpmtc_o,
  output logic              csr_6_o,
  output logic              csr_high_o,

  output logic              mret_o,
  output logic [1:0]        mcause30_o,
  output logic              except_o
);

// This is how custom instructions are smoke-tested. We simply overwrite the
// AND instruction by a custom instruction and implement the AND in the tb ;)
logic [31:0] instr;


//`define SMOKETEST_CCX

`ifdef SMOKETEST_CCX
(* keep *) logic dbg_ccx;
always_comb begin
  if ((instr_i[6:0] == 'b0110011) && (instr_i[14:12] == 'h7)) begin
    instr = {instr_i[21:15], 3'b0, instr_i[11:7], 7'h5B};
  end else begin
    instr = instr_i;
  end
end
assign dbg_ccx = (instr_i != instr);
`else 
assign instr = instr_i;
`endif



// If 1, a smaller decoder is implemented. However, this 
// leads to a reduced fmax
localparam SMALL = 1;

// --- misc ---

logic in_cycle_2;
assign in_cycle_2 = cyc_two_i;

// --- register decoding ---

logic [4:0] rs1_r;
logic [4:0] rs2_r;
logic [4:0] rd_r;

always_ff @(posedge clk_i) begin
  if (~rst_in & (RST != "MIN")) begin
    rs1_r <= 'b0;
    rs2_r <= 'b0;
    rd_r  <= 'b0;
  end else if (stb_ir_i) begin
    rs1_r <= instr[19:15];
    rs2_r <= instr[24:20];
    rd_r  <= instr[11:7];
  end
end

assign rs1_o = rs1_r;
assign rs2_o = rs2_r;
assign rd_o  = rd_r;

assign ccx_sel_o = i_r[13:12];


// --- imm decoding ---

logic [31:0] imm_r, imm_n;

logic [31:0] u_imm;
logic [31:0] j_imm;
logic [31:0] i_imm;
logic [31:0] s_imm;
logic [31:0] b_imm;

assign i_imm = { {21{instr[31]}}, instr[30:20] };
assign s_imm = { {21{instr[31]}}, instr[30:25], instr[11:7] };
assign b_imm = { {20{instr[31]}}, instr[7], instr[30:25],
                  instr[11:8], 1'd0};
assign u_imm = { instr[31:12], 12'd0 };
assign j_imm = { {12{instr[31]}}, instr[19:12], instr[20],
                  instr[30:21], 1'd0 };

logic is_u_imm;
logic is_j_imm;
logic is_i_imm;
logic is_s_imm;
logic is_b_imm;

// TODO: MRET compare are with passthrough + nop in current insn to use
// inc(pc) instead of alu to increment

/* svlint off style_keyword_1or2space */
/* svlint off style_keyword_construct */
/* svlint off style_keyword_1space */
always_comb begin
  imm_n = 32'd4;
  if (is_u_imm) imm_n = u_imm;
  else if (is_j_imm) imm_n = j_imm;
  else if (is_i_imm) imm_n = i_imm;
  else if (is_s_imm) imm_n = s_imm;
  else if (is_b_imm) imm_n = b_imm;
end
/* svlint on style_keyword_1or2space */
/* svlint on style_keyword_construct */
/* svlint on style_keyword_1space */


always_ff @(posedge clk_i) begin
  if (stb_ir_i) begin
    imm_r <= imm_n;
  end else if (shft_imm_i) begin
    imm_r <= {{CHUNKSIZE{1'bx}}, imm_r[31:CHUNKSIZE]};
  end
end

assign imm_o = imm_r[CHUNKSIZE-1:0];

// --- store opcode ---

// let the tool optimize away the bits that are not needed
logic [31:0] i_r;

always_ff @(posedge clk_i) begin
  if (~rst_in) begin
    // either to instr or to NOP, all 0s causes trap
    i_r <= instr; // 'b0;
  end else if (stb_ir_i) begin
    i_r <= instr;
  end
end

// --- masks ---

assign ls_w_o = i_r[13];
assign ls_h_o = i_r[12];
assign ls_b_o = ~ls_w_o & ~ls_h_o;

// Smaller than version below, inspired by SERV
assign ls_mask_o[3] = (adr_lsbs_i == 2'b11) | ls_w_o | (ls_h_o & adr_lsbs_i[1]);
assign ls_mask_o[2] = (adr_lsbs_i == 2'b10) | ls_w_o;
assign ls_mask_o[1] = (adr_lsbs_i == 2'b01) | ls_w_o | (ls_h_o & !adr_lsbs_i[1]);
assign ls_mask_o[0] = (adr_lsbs_i == 2'b00);

//always_comb begin
//  ls_mask_o = 4'b0011;
//  if (ls_w_o) begin
//    ls_mask_o = '1;
//  end else if (ls_h_o) begin
//    if (adr_lsbs_i[1]) begin
//      ls_mask_o = 4'b1100;
//    end
//  end else begin
//    ls_mask_o = (4'b0001 << adr_lsbs_i);
//  end
//end

assign ld_sext_o = i_r[14];
assign sext_o    = (~i_r[14] & ~i_r[4]) | (i_r[30] & i_r[4]);

generate
  if (SMALL) begin
    always_comb begin
      is_b_imm = 1'b0;
      is_s_imm = 1'b0;
      is_i_imm = 1'b0;
      is_j_imm = 1'b0;
      is_u_imm = 1'b0;

      if (instr[2] & instr[3])
        is_j_imm = 1'b1;
      else if (~instr[2] & ~instr[4] & instr[6])
        is_b_imm = 1'b1;
      else if (instr[2] & ~instr[6])
        is_u_imm = 1'b1;
      else if (~instr[2] & ~instr[4] & instr[5])
        is_s_imm = 1'b1;
      // This does not work for csrrxi anymore, but fixes mret efficiently
      //else if (~(instr[4] & instr[5] & ~instr[6]))
      else if (~(instr[4] & instr[5]))
        is_i_imm = 1'b1;

    end
  end else begin

    assign is_b_imm = (!instr[13]&instr[6]&instr[5]&!instr[4]&
        !instr[3]&!instr[2]&instr[1]&instr[0]) | (
        instr[14]&instr[6]&instr[5]&!instr[4]&!instr[3]
        &!instr[2]&instr[1]&instr[0]);

    assign is_s_imm = (!instr[14]&!instr[12]&!instr[6]&instr[5]&
        !instr[4]&!instr[3]&!instr[2]
        &instr[1]&instr[0]) | (!instr[14]&!instr[13]&!instr[6]&
        instr[5]&!instr[4]&!instr[3]
        &!instr[2]&instr[1]&instr[0]);

    assign is_i_imm = (!instr[31]&!instr[30]&!instr[29]&!instr[28]&
    !instr[27]&!instr[26]&!instr[25]&!instr[6]&!instr[5]&instr[4
    ]&!instr[3]&!instr[2]&instr[1]&instr[0]) | (!instr[31]
        &!instr[29]&!instr[28]&!instr[27]&!instr[26]&!instr[25]&
        instr[14]&!instr[6]&!instr[5]
        &instr[4]&!instr[3]&!instr[2]&instr[1]&instr[0]) |
        (!instr[12]&!instr[6]&!instr[5]
        &instr[4]&!instr[3]&!instr[2]&instr[1]&instr[0]) |
        (!instr[14]&!instr[13]&!instr[12]
        &instr[6]&instr[5]&!instr[4]&!instr[3]&instr[2]&
        instr[1]&instr[0]) | (!instr[14]
        &!instr[12]&!instr[6]&!instr[5]&!instr[3]&!instr[2]&
        instr[1]&instr[0]) | (!instr[13]
        &!instr[6]&!instr[5]&!instr[4]&!instr[3]&!instr[2]&
        instr[1]&instr[0]) | (instr[13]
        &!instr[6]&!instr[5]&instr[4]&!instr[3]&!instr[2]&
        instr[1]&instr[0]);

    assign is_j_imm = (instr[6]&instr[5]&!instr[4]&instr[3]&
    instr[2]&instr[1]&instr[0]);

    assign is_u_imm = (!instr[6]&instr[4]&!instr[3]&instr[2]&
    instr[1]&instr[0]);
end
endgenerate

assign alu_aux_b_spm_d_o = (!i_r[14]&!i_r[12]&!i_r[6]&!i_r[5]&!i_r[4]&!i_r[3]
    &!i_r[2]&in_cycle_2) | (!i_r[13]&i_r[12]&!i_r[6]&i_r[4]&!i_r[3]
    &!i_r[2]&in_cycle_2) | (!i_r[13]&!i_r[6]&!i_r[5]&!i_r[4]&!i_r[3]
    &!i_r[2]&in_cycle_2);

assign alu_aux_rs_b_imm_o = (!i_r[13]&!i_r[6]&!i_r[5]&!i_r[3]&!i_r[2]&!in_cycle_2) | (
    i_r[14]&i_r[6]&i_r[5]&!i_r[4]&!i_r[3]&in_cycle_2) | (!i_r[14]&!i_r[13]
    &!i_r[12]&i_r[6]&i_r[5]&i_r[4]&!i_r[3]&!i_r[2]) | (!i_r[13]&i_r[6]
    &i_r[5]&!i_r[4]&!i_r[3]&in_cycle_2) | (i_r[6]&i_r[5]&!i_r[4]&i_r[2]) | (
    !i_r[14]&!i_r[12]&!i_r[6]&!i_r[4]&!i_r[3]&!i_r[2]&!in_cycle_2) | (
    !i_r[14]&!i_r[13]&!i_r[6]&!i_r[4]&!i_r[3]&!i_r[2]&!in_cycle_2) | (
    i_r[13]&!i_r[6]&!i_r[5]&i_r[4]&!i_r[3]) | (!i_r[12]&!i_r[6]&!i_r[5]
    &i_r[4]&!i_r[3]) | (!i_r[6]&i_r[4]&!i_r[3]&i_r[2]);

assign alu_aux_rs_a_pc_o = (!i_r[13]&i_r[6]&i_r[5]&!i_r[4]&!i_r[3]&in_cycle_2) | (
    i_r[14]&i_r[6]&i_r[5]&!i_r[4]&!i_r[3]&in_cycle_2) | (!i_r[6]&i_r[4]
    &!i_r[3]&i_r[2]) | (i_r[6]&i_r[5]&!i_r[4]&i_r[3]&i_r[2]) | (i_r[6]
    &i_r[5]&!i_r[4]&i_r[2]&in_cycle_2) | (trap_entry_i);

assign alu_aux_rev_o = (!i_r[13]&i_r[12]&!i_r[6]&i_r[4]&!i_r[3]&!i_r[2]
    &!in_cycle_2) | (i_r[6]&i_r[5]&!i_r[4]&i_r[2]) | (!i_r[14]&i_r[6]
    &i_r[5]&i_r[4]&!i_r[3]&!i_r[2]&!in_cycle_2) | (trap_entry_i);

assign alu_cmp_inv_o = (!i_r[14]&!i_r[13]&i_r[12]&i_r[5]&!i_r[3]&!i_r[2]) | (
    i_r[14]&i_r[12]&i_r[6]&i_r[5]&!i_r[4]&!i_r[3]);

assign alu_cmp_eq_o = (!i_r[14]&!i_r[13]&i_r[5]&!i_r[3]&!i_r[2]);

assign alu_cmp_sign_o = (!i_r[12]&!i_r[6]&i_r[4]&!i_r[3]) | (!i_r[13]&i_r[6]
    &i_r[5]&!i_r[4]&!i_r[3]);

assign alu_and_o = (!trap_entry_i&i_r[12]&!i_r[6]&i_r[4]&!i_r[3]);

assign alu_xor_o = (!trap_entry_i&!i_r[13]&!i_r[6]&i_r[4]&!i_r[3]);

assign alu_sub_o = (!trap_entry_i&i_r[30]&!i_r[12]&!i_r[6]&i_r[5]&i_r[4]&!i_r[3]
    &!i_r[2]);

assign alu_en_a_o = (!trap_entry_i&!i_r[14]&!i_r[13]&i_r[5]&!i_r[4]&!i_r[3]
    &!i_r[2]&!in_cycle_2) | (!trap_entry_i&!i_r[14]&!i_r[13]&!i_r[12]
    &i_r[5]&i_r[4]&!i_r[3]&!i_r[2]) | (!trap_entry_i&i_r[14]&i_r[6]
    &i_r[5]&!i_r[4]&!i_r[3]&!i_r[2]) | (!trap_entry_i&!i_r[13]&i_r[6]
    &i_r[5]&!i_r[4]&!i_r[3]&!i_r[2]) | (!trap_entry_i&!i_r[13]&!i_r[6]
    &!i_r[5]&!i_r[4]&!i_r[3]&!i_r[2]&!in_cycle_2) | (!trap_entry_i&i_r[6]
    &i_r[5]&!i_r[4]&i_r[2]&!in_cycle_2) | (!trap_entry_i&!i_r[14]&!i_r[12]
    &!i_r[6]&!i_r[3]&!i_r[2]&!in_cycle_2) | (!trap_entry_i&i_r[13]&!i_r[6]
    &i_r[4]&!i_r[3]&!i_r[2]) | (!trap_entry_i&!i_r[12]&!i_r[6]&i_r[4]
    &!i_r[3]&!i_r[2]) | (!trap_entry_i&!i_r[6]&!i_r[5]&i_r[4]&!i_r[3]
    &i_r[2]);

assign alu_arith_o = (!i_r[14]&!i_r[13]&i_r[5]&!i_r[3]&!i_r[2]) | (!i_r[13]
    &i_r[12]&!i_r[6]&i_r[4]&!i_r[3]) | (i_r[14]&i_r[6]&i_r[5]&!i_r[4]
    &!i_r[3]) | (!i_r[14]&i_r[5]&i_r[4]&!i_r[3]&!i_r[2]) | (!i_r[14]
    &!i_r[12]&!i_r[6]&!i_r[3]&!i_r[2]) | (i_r[6]&i_r[5]&!i_r[4]&i_r[2]) | (
    !i_r[13]&!i_r[6]&!i_r[5]&!i_r[4]&!i_r[3]&!i_r[2]) | (!i_r[6]&i_r[4]
    &!i_r[3]&i_r[2]) | (trap_entry_i);

assign instr_jmp_o = (!trap_entry_i&i_r[6]&i_r[5]&!i_r[4]&i_r[2]);

assign instr_any_br_o = (!trap_entry_i&!i_r[13]&i_r[6]&i_r[5]&!i_r[4]&!i_r[3]
    &!i_r[2]) | (!trap_entry_i&i_r[14]&i_r[6]&i_r[5]&!i_r[4]&!i_r[3]
    &!i_r[2]);

assign alu_aux_use_cmp_o = (!trap_entry_i&!i_r[14]&i_r[13]&!i_r[6]&i_r[4]&!i_r[3]
    &!i_r[2]);

assign instr_left_o = (!trap_entry_i&!i_r[14]&!i_r[6]&i_r[4]&!i_r[3]);

assign instr_shft_o = (!trap_entry_i&!i_r[13]&i_r[12]&!i_r[6]&i_r[4]&!i_r[3]
    &!i_r[2]);

assign instr_st_o = (!trap_entry_i&!i_r[14]&!i_r[12]&!i_r[6]&i_r[5]&!i_r[4]
    &!i_r[3]&!i_r[2]) | (!trap_entry_i&!i_r[14]&!i_r[13]&!i_r[6]&i_r[5]
    &!i_r[4]&!i_r[3]&!i_r[2]);

assign instr_ld_o = (!trap_entry_i&!i_r[14]&!i_r[12]&!i_r[6]&!i_r[5]&!i_r[4]
    &!i_r[3]&!i_r[2]) | (!trap_entry_i&!i_r[13]&!i_r[6]&!i_r[5]&!i_r[4]
    &!i_r[3]&!i_r[2]);

assign instr_slt_o = (!trap_entry_i&!i_r[14]&i_r[13]&!i_r[6]&i_r[4]&!i_r[3]
    &!i_r[2]);

assign rf_we_o = (!i_r[6]&i_r[4]&!i_r[3]) | (i_r[6]&i_r[5]&!i_r[4]&i_r[2]) | (
    !i_r[14]&i_r[13]&i_r[5]&i_r[4]&!i_r[3]&!i_r[2]) | (!i_r[14]&!i_r[12]
    &!i_r[6]&!i_r[5]&!i_r[3]&!i_r[2]) | (!i_r[13]&!i_r[6]&!i_r[5]&!i_r[3]
    &!i_r[2]) | (!i_r[14]&i_r[12]&i_r[5]&i_r[4]&!i_r[3]&!i_r[2]) | (
    !i_r[14]&i_r[6]&!i_r[5]&i_r[4]&i_r[3]&!i_r[2]) | (trap_entry_i);

assign ccx_o = (!trap_entry_i&!i_r[14]&i_r[6]&!i_r[5]&i_r[4]&i_r[3]&!i_r[2]);

generate
  if (CONF == "CSR") begin
    assign instr_csr_o = (!trap_entry_i&!i_r[14]&i_r[13]&i_r[6]&i_r[5]&i_r[4]&!i_r[3]
    &!i_r[2]) | (!trap_entry_i&!i_r[14]&i_r[12]&i_r[6]&i_r[5]&i_r[4]
    &!i_r[3]&!i_r[2]);
    assign csr_hpmtc_o  = i_r[31];
    assign csr_6_o      = i_r[26];
    assign csr_high_o   = i_r[27];
  end else begin
    assign instr_csr_o  = 1'b0;
    assign csr_hpmtc_o  = 1'b0;
    assign csr_6_o      = 1'b0;
    assign csr_high_o   = 1'b0;
  end

  if ((CONF == "INT") | (CONF == "CSR")) begin
    assign mret_o = (!trap_entry_i&i_r[29]&!i_r[14]&!i_r[13]&!i_r[12]&i_r[6]&i_r[5]
    &i_r[4]&!i_r[3]&!i_r[2]);
  end else begin
    assign mret_o = 1'b0;
  end
endgenerate

// --- csr and trap ---

generate
  if ((CONF == "CSR") || (CONF == "INT")) begin
    // Illegal instruction: all 0s or all 1s, others might fail to be detected
    // due to area optimization.
    logic trap_insn;
    logic trap_e;

    assign trap_insn  = (&i_r[6:3]) | ~(|i_r[1:0]);
    assign trap_e     = (&i_r[6:4]) &  ~(|i_r[14:12]) & ~i_r[29];
    assign except_o   = trap_insn | trap_e;

    // 2  0010 ... illegal instr
    // 3  0011 ... break
    // 11 1011 ... ecall
    assign mcause30_o[0]  = trap_e;
    assign mcause30_o[1]  = trap_e & i_r[20];

  end else begin
    assign except_o     = 1'b0;
    assign mcause30_o   = 2'b0;
  end
endgenerate


endmodule
